interface myBus (input clk);
  logic [7:0]  data;
  logic      enable;
 
  // From TestBench perspective, 'data' is input and 'write' is output
  // modport TB  (input data, clk, output enable);  
 
  // From DUT perspective, 'data' is output and 'enable' is input
   modport DUT (output data, input enable, clk); 
endinterface


module interface_s (myBus busIf);
  always @ (posedge busIf.clk)
    if (busIf.enable)
      busIf.data <= busIf.data+1;
    else
      busIf.data <= 0;
endmodule


